module draw_grid(values, x, y);
	input [16*4 : 0] values; // all values in order
	output [6:0] x, y; // x: 57-123; y: 27-93.
	
	
endmodule


