module resultdisplay(status);
//TODO: display result and ask to play again
endmodule